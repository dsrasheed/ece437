// interface include
`include "exec_stage_if.vh"

// memory types
`include "cpu_types_pkg.vh"

module exec_stage (
  input CLK, nRST,
  exec_stage.es esif
);

import cpu_types_pkg::*;



endmodule
